module template (
    /*
    input a;
    output reg out;
    */
);

// assign out = a;

endmodule
